library verilog;
use verilog.vl_types.all;
entity MIPS_TB is
end MIPS_TB;
